// Authors : 
//	Harshad Bhausaheb Ugale
//	Mahesh Shahaji Patil

// Description :
//	This module reads memory and gived data.


module Memory_Access
(
	input resetn,flush,
	input [36:0] MemAccessInData,
	
);
